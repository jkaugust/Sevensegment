
`ifndef MONITOR__SV
`define MONITOR__SV


class monitor;
  virtual segintf.TEST vTEST; 
  mailbox mon2scb;
  logic [6:0] outrcv;
  
  function new(mailbox mon2scb,virtual segintf.TEST vTEST); 
     this.vTEST = vTEST; 
     if(mon2scb == null) 
       begin 
         $display(" **ERROR**: mon2scb is null"); 
         $finish; 
       end 
       else 
       this.mon2scb = mon2scb; 
  endfunction : new 
  
  task run();
    forever begin
      wait(vTEST.cr.segout)
      outrcv <= vTEST.cr.segout;
      $display(" %0d : Receiver : Received a segout %0d",$time,outrcv);
      mon2scb.put(outrcv); 
      outrcv <= 7'b0000000; 
    end
   endtask : run
    
endclass : monitor


`endif // MONITOR__SV

