`ifndef DRIVER__SV
`define DRIVER__SV

`include "transactor.sv"

class driver;

  virtual segintf.TEST vTEST; 
  mailbox gen2drv;
  event drv2gen;
  mailbox drv2scb; 
  transactor tr;
  
  function new(input mailbox gen2drv,mailbox drv2scb,input event drv2gen, virtual segintf.TEST vTEST);
  this.gen2drv = gen2drv;
  this.drv2gen=drv2gen;
  this.vTEST = vTEST;
  if(drv2scb == null) 
    begin 
      $display(" **ERROR**: drv2scb is null"); 
      $finish; 
     end 
    else 
  this.drv2scb = drv2scb; 
  endfunction:new
 
  task run();
    forever begin
    gen2drv.peek(tr);
    @(posedge vTEST.clk);
    vTEST.cr.segin <= tr.segin;
    vTEST.cr.en <= tr.en;
    
    drv2scb.put(tr);
    
    gen2drv.get(tr);     // Remove cell from the mailbox
     // ->drv2gen;	   
  end 
    
  endtask :run
 
endclass : driver
`endif // DRIVER__SV


